magic
tech sky130A
magscale 1 2
timestamp 1729214622
<< nwell >>
rect -176 -1500 822 1360
<< nsubdiff >>
rect -140 1290 -78 1324
rect 725 1290 786 1324
rect -140 1261 -106 1290
rect 752 1261 786 1290
rect -140 -1430 -106 -1404
rect 752 -1430 786 -1404
rect -140 -1464 -78 -1430
rect 725 -1464 786 -1430
<< nsubdiffcont >>
rect -78 1290 725 1324
rect -140 -1404 -106 1261
rect 752 -1404 786 1261
rect -78 -1464 725 -1430
<< poly >>
rect -56 1252 36 1268
rect -56 1218 -40 1252
rect -6 1218 36 1252
rect -56 1202 36 1218
rect 6 1174 36 1202
rect 610 1252 702 1268
rect 610 1218 652 1252
rect 686 1218 702 1252
rect 610 1202 702 1218
rect 610 1191 640 1202
rect 94 574 294 674
rect -56 558 36 574
rect -56 524 -40 558
rect -6 524 36 558
rect -56 508 36 524
rect 6 496 36 508
rect 610 558 702 574
rect 610 524 652 558
rect 686 524 702 558
rect 610 508 702 524
rect 610 501 640 508
rect 94 -120 552 -20
rect 6 -648 36 -620
rect -56 -664 36 -648
rect -56 -698 -40 -664
rect -6 -698 36 -664
rect -56 -714 36 -698
rect 610 -648 640 -620
rect 610 -664 702 -648
rect 610 -698 652 -664
rect 686 -698 702 -664
rect 610 -714 702 -698
rect 352 -814 552 -714
rect 6 -1342 36 -1314
rect -56 -1358 36 -1342
rect -56 -1392 -40 -1358
rect -6 -1392 36 -1358
rect -56 -1408 36 -1392
rect 610 -1342 640 -1314
rect 610 -1358 702 -1342
rect 610 -1392 652 -1358
rect 686 -1392 702 -1358
rect 610 -1408 702 -1392
<< polycont >>
rect -40 1218 -6 1252
rect 652 1218 686 1252
rect -40 524 -6 558
rect 652 524 686 558
rect -40 -698 -6 -664
rect 652 -698 686 -664
rect -40 -1392 -6 -1358
rect 652 -1392 686 -1358
<< locali >>
rect -140 1290 -78 1324
rect 725 1290 786 1324
rect -140 1261 -106 1290
rect 752 1261 786 1290
rect -56 1218 -40 1252
rect -6 1218 10 1252
rect 636 1218 652 1252
rect 686 1218 702 1252
rect -40 1174 -6 1218
rect 652 1167 686 1218
rect -56 524 -40 558
rect -6 524 10 558
rect 636 524 652 558
rect 686 524 702 558
rect -40 471 -6 524
rect 652 469 686 524
rect -40 -664 -6 -620
rect 652 -664 686 -620
rect -56 -698 -40 -664
rect -6 -698 10 -664
rect 636 -698 652 -664
rect 686 -698 702 -664
rect -40 -1358 -6 -1314
rect 652 -1358 686 -1314
rect -56 -1392 -40 -1358
rect -6 -1392 10 -1358
rect 636 -1392 652 -1358
rect 686 -1392 702 -1358
rect -140 -1430 -106 -1404
rect 752 -1430 786 -1404
rect -140 -1464 -78 -1430
rect 725 -1464 786 -1430
<< viali >>
rect 652 1290 686 1324
rect -40 1218 -6 1252
rect 652 1218 686 1252
rect -40 524 -6 558
rect 652 524 686 558
rect -40 -698 -6 -664
rect 652 -698 686 -664
rect -40 -1392 -6 -1358
rect 652 -1392 686 -1358
rect -40 -1464 -6 -1430
<< metal1 >>
rect 640 1324 698 1330
rect 640 1290 652 1324
rect 686 1290 698 1324
rect -52 1252 6 1258
rect -52 1218 -40 1252
rect -6 1218 6 1252
rect -52 1212 6 1218
rect 640 1252 698 1290
rect 640 1218 652 1252
rect 686 1218 698 1252
rect 640 1212 698 1218
rect -46 1171 0 1212
rect 646 1174 692 1212
rect -46 1159 88 1171
rect -59 783 -49 1159
rect 3 783 88 1159
rect -46 771 88 783
rect 300 724 345 1171
rect 558 774 692 1174
rect 564 724 598 774
rect 300 690 598 724
rect -52 558 6 564
rect -52 524 -40 558
rect -6 524 6 558
rect -52 518 6 524
rect -46 465 0 518
rect -46 89 39 465
rect 91 89 101 465
rect -46 77 91 89
rect 48 -170 147 -136
rect 48 -217 82 -170
rect -46 -617 88 -217
rect -46 -658 0 -617
rect -52 -664 6 -658
rect -52 -698 -40 -664
rect -6 -698 6 -664
rect -52 -704 6 -698
rect 300 -830 345 690
rect 640 558 698 564
rect 640 524 652 558
rect 686 524 698 558
rect 640 518 698 524
rect 646 477 692 518
rect 558 77 692 477
rect 564 30 598 77
rect 504 -4 598 30
rect 558 -229 692 -217
rect 545 -605 555 -229
rect 607 -605 692 -229
rect 558 -617 692 -605
rect 646 -658 692 -617
rect 640 -664 698 -658
rect 640 -698 652 -664
rect 686 -698 698 -664
rect 640 -704 698 -698
rect 48 -864 345 -830
rect 48 -911 82 -864
rect -46 -1311 88 -911
rect 300 -1311 345 -864
rect 558 -923 692 -911
rect 558 -1299 643 -923
rect 695 -1299 705 -923
rect 558 -1311 692 -1299
rect -46 -1352 0 -1311
rect 646 -1352 692 -1311
rect -52 -1358 6 -1352
rect -52 -1392 -40 -1358
rect -6 -1392 6 -1358
rect -52 -1430 6 -1392
rect 640 -1358 698 -1352
rect 640 -1392 652 -1358
rect 686 -1392 698 -1358
rect 640 -1398 698 -1392
rect -52 -1464 -40 -1430
rect -6 -1464 6 -1430
rect -52 -1470 6 -1464
<< via1 >>
rect -49 783 3 1159
rect 39 89 91 465
rect 555 -605 607 -229
rect 643 -1299 695 -923
<< metal2 >>
rect -49 1159 3 1169
rect -49 665 3 783
rect -53 655 7 665
rect 630 595 639 655
rect 699 595 708 655
rect -53 585 7 595
rect -49 -725 3 585
rect 39 465 91 475
rect 39 -44 91 89
rect 39 -96 607 -44
rect 555 -229 607 -96
rect 555 -615 607 -605
rect 643 -724 695 595
rect -53 -734 7 -725
rect -53 -803 7 -794
rect 639 -734 699 -724
rect 639 -804 699 -794
rect 643 -923 695 -804
rect 643 -1309 695 -1299
<< via2 >>
rect -53 595 7 655
rect 639 595 699 655
rect -53 -794 7 -734
rect 639 -794 699 -734
<< metal3 >>
rect -63 655 17 660
rect 634 655 704 660
rect -63 595 -53 655
rect 7 595 639 655
rect 699 595 704 655
rect -63 590 17 595
rect 634 590 704 595
rect -58 -734 12 -729
rect 629 -734 709 -729
rect -58 -794 -53 -734
rect 7 -794 639 -734
rect 699 -794 709 -734
rect -58 -799 12 -794
rect 629 -799 709 -794
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729133713
transform 1 0 625 0 1 277
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729133713
transform 1 0 21 0 1 -1111
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729133713
transform 1 0 625 0 1 -1111
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729133713
transform 1 0 21 0 1 -417
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729133713
transform 1 0 625 0 1 -417
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729133713
transform 1 0 21 0 1 277
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729133713
transform 1 0 625 0 1 971
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729133713
transform 1 0 21 0 1 971
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729137990
transform 1 0 323 0 1 -1111
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729137990
transform 1 0 323 0 1 -417
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729137990
transform 1 0 323 0 1 277
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729137990
transform 1 0 323 0 1 971
box -323 -300 323 300
<< labels >>
flabel metal2 678 -58 678 -58 0 FreeSans 160 0 0 0 D5
port 0 nsew
flabel metal1 578 16 578 16 0 FreeSans 160 0 0 0 D2
port 1 nsew
flabel metal2 574 -90 574 -90 0 FreeSans 160 0 0 0 D1
port 2 nsew
flabel metal1 670 1276 670 1276 0 FreeSans 160 0 0 0 VDD
port 3 nsew
<< end >>
