magic
tech sky130A
magscale 1 2
timestamp 1729427460
<< psubdiff >>
rect -176 718 -113 752
rect 1046 718 1106 752
rect -176 690 -142 718
rect 1072 690 1106 718
rect -176 -31 -142 4
rect 1072 -31 1106 4
rect -176 -65 -113 -31
rect 1046 -65 1106 -31
<< psubdiffcont >>
rect -113 718 1046 752
rect -176 4 -142 690
rect 1072 4 1106 690
rect -113 -65 1046 -31
<< poly >>
rect -92 671 0 687
rect -92 637 -76 671
rect -42 637 0 671
rect -92 621 0 637
rect -30 618 0 621
rect 930 670 1022 686
rect 930 636 972 670
rect 1006 636 1022 670
rect 930 620 1022 636
rect -92 50 0 66
rect -92 16 -76 50
rect -42 16 0 50
rect -92 0 0 16
rect 930 50 1022 66
rect 930 16 972 50
rect 1006 16 1022 50
rect 930 0 1022 16
<< polycont >>
rect -76 637 -42 671
rect 972 636 1006 670
rect -76 16 -42 50
rect 972 16 1006 50
<< locali >>
rect -176 718 -113 752
rect 1046 718 1106 752
rect -176 690 -142 718
rect 1072 690 1106 718
rect -92 637 -76 671
rect -42 637 -26 671
rect 956 636 972 670
rect 1006 636 1022 670
rect -92 16 -76 50
rect -42 16 -26 50
rect 956 16 972 50
rect 1006 16 1022 50
rect -176 -31 -142 4
rect 1072 -31 1106 4
rect -176 -65 -113 -31
rect 1046 -65 1106 -31
<< viali >>
rect 230 718 264 752
rect 666 718 700 752
rect -76 637 -42 671
rect 972 636 1006 670
rect -76 16 -42 50
rect 972 16 1006 50
rect 230 -65 264 -31
rect 666 -65 700 -31
<< metal1 >>
rect 218 752 276 758
rect 218 718 230 752
rect 264 718 276 752
rect 218 712 276 718
rect 654 752 712 758
rect 654 718 666 752
rect 700 718 712 752
rect 654 712 712 718
rect -88 671 -30 677
rect -88 637 -76 671
rect -42 637 -30 671
rect -88 631 -30 637
rect -82 598 -36 631
rect -82 398 52 598
rect 230 582 264 712
rect 429 410 439 586
rect 491 410 501 586
rect 666 582 700 712
rect 960 670 1018 676
rect 960 636 972 670
rect 1006 636 1018 670
rect 960 630 1018 636
rect 966 598 1012 630
rect 6 366 52 398
rect 878 398 1012 598
rect 878 366 924 398
rect 6 320 86 366
rect 162 320 777 365
rect 845 320 924 366
rect -82 276 52 288
rect -82 100 3 276
rect 55 100 65 276
rect 442 273 487 320
rect 878 276 1012 288
rect -82 88 52 100
rect -82 56 -36 88
rect -88 50 -30 56
rect -88 16 -76 50
rect -42 16 -30 50
rect -88 10 -30 16
rect 230 -25 264 110
rect 865 100 875 276
rect 927 100 1012 276
rect 666 -25 700 91
rect 878 88 1012 100
rect 966 56 1012 88
rect 960 50 1018 56
rect 960 16 972 50
rect 1006 16 1018 50
rect 960 10 1018 16
rect 218 -31 276 -25
rect 218 -65 230 -31
rect 264 -65 276 -31
rect 218 -71 276 -65
rect 654 -31 712 -25
rect 654 -65 666 -31
rect 700 -65 712 -31
rect 654 -71 712 -65
<< via1 >>
rect 439 410 491 586
rect 3 100 55 276
rect 875 100 927 276
<< metal2 >>
rect 439 586 491 596
rect 439 369 491 410
rect 3 317 927 369
rect 3 276 55 317
rect 3 90 55 100
rect 875 276 927 317
rect 875 90 927 100
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1729427460
transform 1 0 -15 0 1 498
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729427460
transform 1 0 945 0 1 498
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729427460
transform 1 0 945 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729427460
transform 1 0 -15 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_YYNGNX  sky130_fd_pr__nfet_01v8_YYNGNX_0
timestamp 1729427460
transform 1 0 465 0 1 343
box -465 -343 465 343
<< labels >>
flabel metal1 27 386 27 386 0 FreeSans 1600 0 0 0 D8
port 1 nsew
flabel metal2 900 300 900 300 0 FreeSans 1600 0 0 0 D9
port 2 nsew
flabel metal1 682 -3 682 -3 0 FreeSans 480 0 0 0 gnd
port 3 nsew
<< end >>
