magic
tech sky130A
magscale 1 2
timestamp 1729427460
<< nmos >>
rect -407 55 -247 255
rect -189 55 -29 255
rect 29 55 189 255
rect 247 55 407 255
rect -407 -255 -247 -55
rect -189 -255 -29 -55
rect 29 -255 189 -55
rect 247 -255 407 -55
<< ndiff >>
rect -465 243 -407 255
rect -465 67 -453 243
rect -419 67 -407 243
rect -465 55 -407 67
rect -247 243 -189 255
rect -247 67 -235 243
rect -201 67 -189 243
rect -247 55 -189 67
rect -29 243 29 255
rect -29 67 -17 243
rect 17 67 29 243
rect -29 55 29 67
rect 189 243 247 255
rect 189 67 201 243
rect 235 67 247 243
rect 189 55 247 67
rect 407 243 465 255
rect 407 67 419 243
rect 453 67 465 243
rect 407 55 465 67
rect -465 -67 -407 -55
rect -465 -243 -453 -67
rect -419 -243 -407 -67
rect -465 -255 -407 -243
rect -247 -67 -189 -55
rect -247 -243 -235 -67
rect -201 -243 -189 -67
rect -247 -255 -189 -243
rect -29 -67 29 -55
rect -29 -243 -17 -67
rect 17 -243 29 -67
rect -29 -255 29 -243
rect 189 -67 247 -55
rect 189 -243 201 -67
rect 235 -243 247 -67
rect 189 -255 247 -243
rect 407 -67 465 -55
rect 407 -243 419 -67
rect 453 -243 465 -67
rect 407 -255 465 -243
<< ndiffc >>
rect -453 67 -419 243
rect -235 67 -201 243
rect -17 67 17 243
rect 201 67 235 243
rect 419 67 453 243
rect -453 -243 -419 -67
rect -235 -243 -201 -67
rect -17 -243 17 -67
rect 201 -243 235 -67
rect 419 -243 453 -67
<< poly >>
rect -407 327 -247 343
rect -407 293 -391 327
rect -263 293 -247 327
rect -407 255 -247 293
rect -189 327 -29 343
rect -189 293 -173 327
rect -45 293 -29 327
rect -189 255 -29 293
rect 29 327 189 343
rect 29 293 45 327
rect 173 293 189 327
rect 29 255 189 293
rect 247 327 407 343
rect 247 293 263 327
rect 391 293 407 327
rect 247 255 407 293
rect -407 17 -247 55
rect -407 -17 -391 17
rect -263 -17 -247 17
rect -407 -55 -247 -17
rect -189 17 -29 55
rect -189 -17 -173 17
rect -45 -17 -29 17
rect -189 -55 -29 -17
rect 29 17 189 55
rect 29 -17 45 17
rect 173 -17 189 17
rect 29 -55 189 -17
rect 247 17 407 55
rect 247 -17 263 17
rect 391 -17 407 17
rect 247 -55 407 -17
rect -407 -293 -247 -255
rect -407 -327 -391 -293
rect -263 -327 -247 -293
rect -407 -343 -247 -327
rect -189 -293 -29 -255
rect -189 -327 -173 -293
rect -45 -327 -29 -293
rect -189 -343 -29 -327
rect 29 -293 189 -255
rect 29 -327 45 -293
rect 173 -327 189 -293
rect 29 -343 189 -327
rect 247 -293 407 -255
rect 247 -327 263 -293
rect 391 -327 407 -293
rect 247 -343 407 -327
<< polycont >>
rect -391 293 -263 327
rect -173 293 -45 327
rect 45 293 173 327
rect 263 293 391 327
rect -391 -17 -263 17
rect -173 -17 -45 17
rect 45 -17 173 17
rect 263 -17 391 17
rect -391 -327 -263 -293
rect -173 -327 -45 -293
rect 45 -327 173 -293
rect 263 -327 391 -293
<< locali >>
rect -407 293 -391 327
rect -263 293 -247 327
rect -189 293 -173 327
rect -45 293 -29 327
rect 29 293 45 327
rect 173 293 189 327
rect 247 293 263 327
rect 391 293 407 327
rect -453 243 -419 259
rect -453 51 -419 67
rect -235 243 -201 259
rect -235 51 -201 67
rect -17 243 17 259
rect -17 51 17 67
rect 201 243 235 259
rect 201 51 235 67
rect 419 243 453 259
rect 419 51 453 67
rect -407 -17 -391 17
rect -263 -17 -247 17
rect -189 -17 -173 17
rect -45 -17 -29 17
rect 29 -17 45 17
rect 173 -17 189 17
rect 247 -17 263 17
rect 391 -17 407 17
rect -453 -67 -419 -51
rect -453 -259 -419 -243
rect -235 -67 -201 -51
rect -235 -259 -201 -243
rect -17 -67 17 -51
rect -17 -259 17 -243
rect 201 -67 235 -51
rect 201 -259 235 -243
rect 419 -67 453 -51
rect 419 -259 453 -243
rect -407 -327 -391 -293
rect -263 -327 -247 -293
rect -189 -327 -173 -293
rect -45 -327 -29 -293
rect 29 -327 45 -293
rect 173 -327 189 -293
rect 247 -327 263 -293
rect 391 -327 407 -293
<< viali >>
rect -372 293 -282 327
rect -154 293 -64 327
rect 64 293 154 327
rect 282 293 372 327
rect -453 67 -419 243
rect -235 67 -201 243
rect -17 67 17 243
rect 201 67 235 243
rect 419 67 453 243
rect -372 -17 -282 17
rect -154 -17 -64 17
rect 64 -17 154 17
rect 282 -17 372 17
rect -453 -243 -419 -67
rect -235 -243 -201 -67
rect -17 -243 17 -67
rect 201 -243 235 -67
rect 419 -243 453 -67
rect -372 -327 -282 -293
rect -154 -327 -64 -293
rect 64 -327 154 -293
rect 282 -327 372 -293
<< metal1 >>
rect -384 327 -270 333
rect -384 293 -372 327
rect -282 293 -270 327
rect -384 287 -270 293
rect -166 327 -52 333
rect -166 293 -154 327
rect -64 293 -52 327
rect -166 287 -52 293
rect 52 327 166 333
rect 52 293 64 327
rect 154 293 166 327
rect 52 287 166 293
rect 270 327 384 333
rect 270 293 282 327
rect 372 293 384 327
rect 270 287 384 293
rect -459 243 -413 255
rect -459 67 -453 243
rect -419 67 -413 243
rect -459 55 -413 67
rect -241 243 -195 255
rect -241 67 -235 243
rect -201 67 -195 243
rect -241 55 -195 67
rect -23 243 23 255
rect -23 67 -17 243
rect 17 67 23 243
rect -23 55 23 67
rect 195 243 241 255
rect 195 67 201 243
rect 235 67 241 243
rect 195 55 241 67
rect 413 243 459 255
rect 413 67 419 243
rect 453 67 459 243
rect 413 55 459 67
rect -384 17 -270 23
rect -384 -17 -372 17
rect -282 -17 -270 17
rect -384 -23 -270 -17
rect -166 17 -52 23
rect -166 -17 -154 17
rect -64 -17 -52 17
rect -166 -23 -52 -17
rect 52 17 166 23
rect 52 -17 64 17
rect 154 -17 166 17
rect 52 -23 166 -17
rect 270 17 384 23
rect 270 -17 282 17
rect 372 -17 384 17
rect 270 -23 384 -17
rect -459 -67 -413 -55
rect -459 -243 -453 -67
rect -419 -243 -413 -67
rect -459 -255 -413 -243
rect -241 -67 -195 -55
rect -241 -243 -235 -67
rect -201 -243 -195 -67
rect -241 -255 -195 -243
rect -23 -67 23 -55
rect -23 -243 -17 -67
rect 17 -243 23 -67
rect -23 -255 23 -243
rect 195 -67 241 -55
rect 195 -243 201 -67
rect 235 -243 241 -67
rect 195 -255 241 -243
rect 413 -67 459 -55
rect 413 -243 419 -67
rect 453 -243 459 -67
rect 413 -255 459 -243
rect -384 -293 -270 -287
rect -384 -327 -372 -293
rect -282 -327 -270 -293
rect -384 -333 -270 -327
rect -166 -293 -52 -287
rect -166 -327 -154 -293
rect -64 -327 -52 -293
rect -166 -333 -52 -327
rect 52 -293 166 -287
rect 52 -327 64 -293
rect 154 -327 166 -293
rect 52 -333 166 -327
rect 270 -293 384 -287
rect 270 -327 282 -293
rect 372 -327 384 -293
rect 270 -333 384 -327
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 2 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 1 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
