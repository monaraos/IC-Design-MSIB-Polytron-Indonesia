magic
tech sky130A
magscale 1 2
timestamp 1729428309
<< nwell >>
rect 116 3260 2307 3264
rect 0 1932 2770 3260
rect 0 -421 1002 3
<< viali >>
rect 1587 1752 1621 1786
rect 1118 1555 1298 1690
rect 1121 1347 1301 1482
rect 1123 938 1303 1073
rect 1124 506 1304 641
<< metal1 >>
rect 812 3088 872 3094
rect 872 3028 1175 3088
rect 812 3022 872 3028
rect 816 2814 1042 2872
rect 816 2812 874 2814
rect 984 1647 1042 2814
rect 1115 2628 1175 3028
rect 1115 2568 1647 2628
rect 1579 2044 1631 2050
rect 1151 1696 1224 2006
rect 1579 1986 1631 1992
rect 2637 1949 2691 2041
rect 1369 1901 2691 1949
rect 1106 1690 1310 1696
rect 1106 1647 1118 1690
rect 984 1589 1118 1647
rect 1106 1555 1118 1589
rect 1298 1555 1310 1690
rect 1106 1549 1310 1555
rect 691 1496 1053 1530
rect 1019 -6 1053 1496
rect 1109 1482 1313 1488
rect 1109 1347 1121 1482
rect 1301 1444 1313 1482
rect 1369 1444 1423 1901
rect 1656 1525 1666 1701
rect 1718 1525 1728 1701
rect 1301 1390 1423 1444
rect 1301 1347 1313 1390
rect 1109 1341 1313 1347
rect 1113 1140 1123 1275
rect 1303 1140 1313 1275
rect 1111 1073 1315 1082
rect 1111 938 1123 1073
rect 1303 1031 1315 1073
rect 1881 1031 1939 1057
rect 1303 980 2067 1031
rect 1303 938 1315 980
rect 2009 948 2067 980
rect 1111 928 1315 938
rect 1113 723 1123 858
rect 1303 723 1313 858
rect 1112 641 1316 647
rect 1112 506 1124 641
rect 1304 506 1316 641
rect 1112 500 1316 506
rect 1189 306 1245 500
rect 1368 338 1825 371
rect 1183 250 1189 306
rect 1245 250 1251 306
rect 1189 244 1245 250
rect 1368 161 1401 338
rect 1359 155 1411 161
rect 1359 97 1411 103
rect 1264 -6 1270 3
rect 1019 -40 1270 -6
rect 1264 -49 1270 -40
rect 1322 -49 1328 3
<< via1 >>
rect 812 3028 872 3088
rect 1579 1992 1631 2044
rect 1666 1525 1718 1701
rect 1123 1140 1303 1275
rect 1123 723 1303 858
rect 1189 250 1245 306
rect 1359 103 1411 155
rect 1270 -49 1322 3
<< metal2 >>
rect 984 3127 1168 3181
rect 806 3086 812 3088
rect 872 3086 878 3088
rect 805 3030 812 3086
rect 872 3030 879 3086
rect 806 3028 812 3030
rect 872 3028 878 3030
rect 728 1271 784 1281
rect 984 1236 1038 3127
rect 1886 2440 1942 2450
rect 1886 2255 1942 2265
rect 1566 1988 1575 2048
rect 1635 1988 1644 2048
rect 1579 1948 1631 1988
rect 1579 1896 1718 1948
rect 1666 1701 1718 1896
rect 1666 1515 1718 1525
rect 1664 1391 1720 1401
rect 1123 1275 1303 1285
rect 984 1182 1123 1236
rect 1664 1205 1720 1215
rect 1123 1130 1303 1140
rect 728 885 784 895
rect 1123 858 1303 868
rect 1303 765 1406 808
rect 1123 713 1303 723
rect 1187 308 1247 317
rect 1183 250 1187 306
rect 1247 250 1251 306
rect 1363 291 1406 765
rect 1363 248 2042 291
rect 1187 239 1247 248
rect 1346 99 1355 159
rect 1415 99 1424 159
rect 1270 7 1322 9
rect 1257 -53 1266 7
rect 1326 -53 1335 7
rect 1270 -55 1322 -53
<< via2 >>
rect 814 3030 870 3086
rect 728 895 784 1271
rect 1886 2265 1942 2440
rect 1575 2044 1635 2048
rect 1575 1992 1579 2044
rect 1579 1992 1631 2044
rect 1631 1992 1635 2044
rect 1575 1988 1635 1992
rect 1664 1215 1720 1391
rect 1187 306 1247 308
rect 1187 250 1189 306
rect 1189 250 1245 306
rect 1245 250 1247 306
rect 1187 248 1247 250
rect 1355 155 1415 159
rect 1355 103 1359 155
rect 1359 103 1411 155
rect 1411 103 1415 155
rect 1355 99 1415 103
rect 1266 3 1326 7
rect 1266 -49 1270 3
rect 1270 -49 1322 3
rect 1322 -49 1326 3
rect 1266 -53 1326 -49
<< metal3 >>
rect 809 3086 875 3091
rect 809 3030 814 3086
rect 870 3030 875 3086
rect 809 3025 875 3030
rect 812 2951 872 3025
rect 812 2891 1046 2951
rect 986 2155 1046 2891
rect 1876 2440 1952 2445
rect 750 2095 1046 2155
rect 724 1394 1084 1454
rect 724 1276 784 1394
rect 718 1271 794 1276
rect 718 895 728 1271
rect 784 895 794 1271
rect 718 890 794 895
rect 1024 159 1084 1394
rect 1355 1035 1415 2340
rect 1876 2265 1886 2440
rect 1942 2265 1952 2440
rect 1876 2260 1952 2265
rect 1570 2048 1640 2053
rect 1884 2048 1944 2260
rect 1570 1988 1575 2048
rect 1635 1988 1944 2048
rect 1570 1983 1640 1988
rect 1654 1391 1730 1396
rect 1654 1215 1664 1391
rect 1720 1215 1730 1391
rect 1654 1210 1730 1215
rect 1663 1035 1723 1210
rect 1355 975 1723 1035
rect 1182 308 1252 313
rect 1355 308 1415 975
rect 1182 248 1187 308
rect 1247 248 1415 308
rect 1182 243 1252 248
rect 1350 159 1420 164
rect 1024 99 1355 159
rect 1415 99 1420 159
rect 1350 94 1420 99
rect 1261 7 1331 12
rect 1261 -53 1266 7
rect 1326 -53 1513 7
rect 1261 -58 1331 -53
rect 1453 -360 1513 -53
rect 1750 -360 1810 -230
rect 1453 -420 1810 -360
use nmos_diff  nmos_diff_0
timestamp 1729427460
transform 1 0 1663 0 1 1115
box -176 -71 1106 758
use nmoscs  nmoscs_0
timestamp 1729226415
transform 1 0 1751 0 1 321
box -288 -741 1014 647
use pmos_diff  pmos_diff_0
timestamp 1729420276
transform 1 0 1755 0 1 2170
box -721 -232 1016 1091
use pmoscs  pmoscs_0
timestamp 1729214622
transform 1 0 176 0 1 1500
box -176 -1500 822 1360
<< labels >>
flabel viali 1211 1611 1211 1611 0 FreeSans 800 0 0 0 vdd
port 1 nsew
flabel viali 1209 1413 1209 1413 0 FreeSans 800 0 0 0 vin
port 2 nsew
flabel via1 1209 1209 1209 1209 0 FreeSans 800 0 0 0 vip
port 3 nsew
flabel viali 1209 1010 1209 1010 0 FreeSans 800 0 0 0 gnd
port 4 nsew
flabel via1 1213 795 1213 795 0 FreeSans 800 0 0 0 RS
port 5 nsew
flabel viali 1215 568 1215 568 0 FreeSans 800 0 0 0 out
port 6 nsew
<< end >>
